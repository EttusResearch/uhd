//
// Copyright 2021 Ettus Research, a National Instruments Brand
//
// SPDX-License-Identifier: LGPL-3.0-or-later
//
// Module: x4xx_mgt_type.vh
// Description:  Enumerations for types of MGT to be used with the X4XX
//

`define MGT_100GbE       5
`define MGT_WhiteRabbit  4
`define MGT_Aurora       3
`define MGT_10GbE        2
`define MGT_1GbE         1
`define MGT_Disabled     0
