//
// Copyright 2011 Ettus Research LLC
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.
//


// Skeleton PHY interface simulator

module miim_model(input mdc_i, 
		  inout mdio, 
		  input phy_resetn_i, 
		  input phy_clk_i, 
		  output phy_intn_o,
		  output [2:0] speed_o);

   assign 		       phy_intn_o = 1;    // No interrupts
   assign 		       speed_o = 3'b100;  // 1G mode
   
endmodule // miim_model
