
module gpif_rd
  ();
   
endmodule // gpif_rd
