//
// Copyright 2011 Ettus Research LLC
//
// This program is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.
//



module gray2bin
  #(parameter WIDTH=8)
    (input [WIDTH-1:0] gray,
     output reg [WIDTH-1:0] bin);

   integer 		i;
   always @(gray)
     for(i = 0;i<WIDTH;i=i+1)
	  bin[i] = ^(gray>>i);
   
endmodule // gray2bin
