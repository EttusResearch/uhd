//
// Copyright 2024 Ettus Research, a National Instruments Brand
//
// SPDX-License-Identifier: LGPL-3.0-or-later
//
// Package: ctrlport_pkg
//
// Description:
//
//   Defines constants for the control-port interface.
//

package ctrlport_pkg;

  `include "ctrlport.vh"

endpackage : ctrlport_pkg
