//
// Copyright 2024 Ettus Research, a National Instruments Brand
//
// SPDX-License-Identifier: LGPL-3.0-or-later
//
// Module: rfnoc_chdr_utils_pkg
//
// Description:
//
//   Package containing constants and functions for working with CHDR.
//

package rfnoc_chdr_utils_pkg;

  `include "rfnoc_chdr_utils.vh"

endpackage : rfnoc_chdr_utils_pkg
